module PC_LUT #(parameter D=12)(
  input       [4:0] addr,	   // target 4 values
  output logic[D-1:0] target);

  always_comb case(addr)
		
			// Program 1
			1: target = 9;
			2: target = 15;
			3: target = 48;
			4: target = 55;
			5: target = 58;
			6: target = 65;
			7: target = 68;
			8: target = 75;
			9: target = 79;
			10: target = 81;
			11: target = 85;
			12: target = 87;
			13: target = 92;
			14: target = 96;

			// Program 2
			15: target = 14;
			16: target = 30;
			17: target = 52;
			18: target = 57;
			19: target = 75;
			20: target = 65;
			21: target = 70;
			22: target = 86;
			23: target = 95;
			24: target = 121;
			25: target = 124;
			26: target = 138;
			27: target = 146;
			28: target = 160;
			29: target = 168;
			30: target = 172;
			31: target = 176;
	default: target = 'b0;  // hold PC  
  endcase

endmodule